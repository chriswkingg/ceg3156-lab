LIBRARY ieee;
USE  ieee.std_logic_1164.all;

ENTITY ControlUnit is
    PORT
    (

    );
    END ControlUnit;

ARCHITECTURE rtl of ControlUnit is
BEGIN

END ARCHITECTURE;